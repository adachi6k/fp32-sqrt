function logic [15:0] lut_inv_sqrt(input logic [7:0] index);
    case (index)
        8'h00: lut_inv_sqrt = 16'h8000;
        8'h01: lut_inv_sqrt = 16'h7FC0;
        8'h02: lut_inv_sqrt = 16'h7F80;
        8'h03: lut_inv_sqrt = 16'h7F41;
        8'h04: lut_inv_sqrt = 16'h7F02;
        8'h05: lut_inv_sqrt = 16'h7EC4;
        8'h06: lut_inv_sqrt = 16'h7E86;
        8'h07: lut_inv_sqrt = 16'h7E48;
        8'h08: lut_inv_sqrt = 16'h7E0B;
        8'h09: lut_inv_sqrt = 16'h7DCE;
        8'h0A: lut_inv_sqrt = 16'h7D92;
        8'h0B: lut_inv_sqrt = 16'h7D55;
        8'h0C: lut_inv_sqrt = 16'h7D19;
        8'h0D: lut_inv_sqrt = 16'h7CDE;
        8'h0E: lut_inv_sqrt = 16'h7CA3;
        8'h0F: lut_inv_sqrt = 16'h7C68;
        8'h10: lut_inv_sqrt = 16'h7C2D;
        8'h11: lut_inv_sqrt = 16'h7BF3;
        8'h12: lut_inv_sqrt = 16'h7BB9;
        8'h13: lut_inv_sqrt = 16'h7B7F;
        8'h14: lut_inv_sqrt = 16'h7B46;
        8'h15: lut_inv_sqrt = 16'h7B0D;
        8'h16: lut_inv_sqrt = 16'h7AD4;
        8'h17: lut_inv_sqrt = 16'h7A9C;
        8'h18: lut_inv_sqrt = 16'h7A64;
        8'h19: lut_inv_sqrt = 16'h7A2C;
        8'h1A: lut_inv_sqrt = 16'h79F4;
        8'h1B: lut_inv_sqrt = 16'h79BD;
        8'h1C: lut_inv_sqrt = 16'h7986;
        8'h1D: lut_inv_sqrt = 16'h7950;
        8'h1E: lut_inv_sqrt = 16'h7919;
        8'h1F: lut_inv_sqrt = 16'h78E3;
        8'h20: lut_inv_sqrt = 16'h78AD;
        8'h21: lut_inv_sqrt = 16'h7878;
        8'h22: lut_inv_sqrt = 16'h7843;
        8'h23: lut_inv_sqrt = 16'h780E;
        8'h24: lut_inv_sqrt = 16'h77D9;
        8'h25: lut_inv_sqrt = 16'h77A5;
        8'h26: lut_inv_sqrt = 16'h7771;
        8'h27: lut_inv_sqrt = 16'h773D;
        8'h28: lut_inv_sqrt = 16'h7709;
        8'h29: lut_inv_sqrt = 16'h76D6;
        8'h2A: lut_inv_sqrt = 16'h76A3;
        8'h2B: lut_inv_sqrt = 16'h7670;
        8'h2C: lut_inv_sqrt = 16'h763D;
        8'h2D: lut_inv_sqrt = 16'h760B;
        8'h2E: lut_inv_sqrt = 16'h75D9;
        8'h2F: lut_inv_sqrt = 16'h75A7;
        8'h30: lut_inv_sqrt = 16'h7575;
        8'h31: lut_inv_sqrt = 16'h7544;
        8'h32: lut_inv_sqrt = 16'h7513;
        8'h33: lut_inv_sqrt = 16'h74E2;
        8'h34: lut_inv_sqrt = 16'h74B2;
        8'h35: lut_inv_sqrt = 16'h7481;
        8'h36: lut_inv_sqrt = 16'h7451;
        8'h37: lut_inv_sqrt = 16'h7421;
        8'h38: lut_inv_sqrt = 16'h73F1;
        8'h39: lut_inv_sqrt = 16'h73C2;
        8'h3A: lut_inv_sqrt = 16'h7393;
        8'h3B: lut_inv_sqrt = 16'h7364;
        8'h3C: lut_inv_sqrt = 16'h7335;
        8'h3D: lut_inv_sqrt = 16'h7306;
        8'h3E: lut_inv_sqrt = 16'h72D8;
        8'h3F: lut_inv_sqrt = 16'h72AA;
        8'h40: lut_inv_sqrt = 16'h727C;
        8'h41: lut_inv_sqrt = 16'h724E;
        8'h42: lut_inv_sqrt = 16'h7221;
        8'h43: lut_inv_sqrt = 16'h71F4;
        8'h44: lut_inv_sqrt = 16'h71C7;
        8'h45: lut_inv_sqrt = 16'h719A;
        8'h46: lut_inv_sqrt = 16'h716D;
        8'h47: lut_inv_sqrt = 16'h7141;
        8'h48: lut_inv_sqrt = 16'h7114;
        8'h49: lut_inv_sqrt = 16'h70E8;
        8'h4A: lut_inv_sqrt = 16'h70BD;
        8'h4B: lut_inv_sqrt = 16'h7091;
        8'h4C: lut_inv_sqrt = 16'h7066;
        8'h4D: lut_inv_sqrt = 16'h703A;
        8'h4E: lut_inv_sqrt = 16'h700F;
        8'h4F: lut_inv_sqrt = 16'h6FE4;
        8'h50: lut_inv_sqrt = 16'h6FBA;
        8'h51: lut_inv_sqrt = 16'h6F8F;
        8'h52: lut_inv_sqrt = 16'h6F65;
        8'h53: lut_inv_sqrt = 16'h6F3B;
        8'h54: lut_inv_sqrt = 16'h6F11;
        8'h55: lut_inv_sqrt = 16'h6EE7;
        8'h56: lut_inv_sqrt = 16'h6EBE;
        8'h57: lut_inv_sqrt = 16'h6E94;
        8'h58: lut_inv_sqrt = 16'h6E6B;
        8'h59: lut_inv_sqrt = 16'h6E42;
        8'h5A: lut_inv_sqrt = 16'h6E19;
        8'h5B: lut_inv_sqrt = 16'h6DF1;
        8'h5C: lut_inv_sqrt = 16'h6DC8;
        8'h5D: lut_inv_sqrt = 16'h6DA0;
        8'h5E: lut_inv_sqrt = 16'h6D78;
        8'h5F: lut_inv_sqrt = 16'h6D50;
        8'h60: lut_inv_sqrt = 16'h6D28;
        8'h61: lut_inv_sqrt = 16'h6D01;
        8'h62: lut_inv_sqrt = 16'h6CD9;
        8'h63: lut_inv_sqrt = 16'h6CB2;
        8'h64: lut_inv_sqrt = 16'h6C8B;
        8'h65: lut_inv_sqrt = 16'h6C64;
        8'h66: lut_inv_sqrt = 16'h6C3D;
        8'h67: lut_inv_sqrt = 16'h6C16;
        8'h68: lut_inv_sqrt = 16'h6BF0;
        8'h69: lut_inv_sqrt = 16'h6BCA;
        8'h6A: lut_inv_sqrt = 16'h6BA3;
        8'h6B: lut_inv_sqrt = 16'h6B7D;
        8'h6C: lut_inv_sqrt = 16'h6B58;
        8'h6D: lut_inv_sqrt = 16'h6B32;
        8'h6E: lut_inv_sqrt = 16'h6B0C;
        8'h6F: lut_inv_sqrt = 16'h6AE7;
        8'h70: lut_inv_sqrt = 16'h6AC2;
        8'h71: lut_inv_sqrt = 16'h6A9D;
        8'h72: lut_inv_sqrt = 16'h6A78;
        8'h73: lut_inv_sqrt = 16'h6A53;
        8'h74: lut_inv_sqrt = 16'h6A2F;
        8'h75: lut_inv_sqrt = 16'h6A0A;
        8'h76: lut_inv_sqrt = 16'h69E6;
        8'h77: lut_inv_sqrt = 16'h69C2;
        8'h78: lut_inv_sqrt = 16'h699E;
        8'h79: lut_inv_sqrt = 16'h697A;
        8'h7A: lut_inv_sqrt = 16'h6956;
        8'h7B: lut_inv_sqrt = 16'h6932;
        8'h7C: lut_inv_sqrt = 16'h690F;
        8'h7D: lut_inv_sqrt = 16'h68EC;
        8'h7E: lut_inv_sqrt = 16'h68C8;
        8'h7F: lut_inv_sqrt = 16'h68A5;
        8'h80: lut_inv_sqrt = 16'h6882;
        8'h81: lut_inv_sqrt = 16'h6860;
        8'h82: lut_inv_sqrt = 16'h683D;
        8'h83: lut_inv_sqrt = 16'h681B;
        8'h84: lut_inv_sqrt = 16'h67F8;
        8'h85: lut_inv_sqrt = 16'h67D6;
        8'h86: lut_inv_sqrt = 16'h67B4;
        8'h87: lut_inv_sqrt = 16'h6792;
        8'h88: lut_inv_sqrt = 16'h6770;
        8'h89: lut_inv_sqrt = 16'h674E;
        8'h8A: lut_inv_sqrt = 16'h672D;
        8'h8B: lut_inv_sqrt = 16'h670B;
        8'h8C: lut_inv_sqrt = 16'h66EA;
        8'h8D: lut_inv_sqrt = 16'h66C9;
        8'h8E: lut_inv_sqrt = 16'h66A8;
        8'h8F: lut_inv_sqrt = 16'h6687;
        8'h90: lut_inv_sqrt = 16'h6666;
        8'h91: lut_inv_sqrt = 16'h6645;
        8'h92: lut_inv_sqrt = 16'h6625;
        8'h93: lut_inv_sqrt = 16'h6604;
        8'h94: lut_inv_sqrt = 16'h65E4;
        8'h95: lut_inv_sqrt = 16'h65C4;
        8'h96: lut_inv_sqrt = 16'h65A3;
        8'h97: lut_inv_sqrt = 16'h6583;
        8'h98: lut_inv_sqrt = 16'h6564;
        8'h99: lut_inv_sqrt = 16'h6544;
        8'h9A: lut_inv_sqrt = 16'h6524;
        8'h9B: lut_inv_sqrt = 16'h6505;
        8'h9C: lut_inv_sqrt = 16'h64E5;
        8'h9D: lut_inv_sqrt = 16'h64C6;
        8'h9E: lut_inv_sqrt = 16'h64A7;
        8'h9F: lut_inv_sqrt = 16'h6488;
        8'hA0: lut_inv_sqrt = 16'h6469;
        8'hA1: lut_inv_sqrt = 16'h644A;
        8'hA2: lut_inv_sqrt = 16'h642B;
        8'hA3: lut_inv_sqrt = 16'h640D;
        8'hA4: lut_inv_sqrt = 16'h63EE;
        8'hA5: lut_inv_sqrt = 16'h63D0;
        8'hA6: lut_inv_sqrt = 16'h63B1;
        8'hA7: lut_inv_sqrt = 16'h6393;
        8'hA8: lut_inv_sqrt = 16'h6375;
        8'hA9: lut_inv_sqrt = 16'h6357;
        8'hAA: lut_inv_sqrt = 16'h6339;
        8'hAB: lut_inv_sqrt = 16'h631C;
        8'hAC: lut_inv_sqrt = 16'h62FE;
        8'hAD: lut_inv_sqrt = 16'h62E0;
        8'hAE: lut_inv_sqrt = 16'h62C3;
        8'hAF: lut_inv_sqrt = 16'h62A6;
        8'hB0: lut_inv_sqrt = 16'h6288;
        8'hB1: lut_inv_sqrt = 16'h626B;
        8'hB2: lut_inv_sqrt = 16'h624E;
        8'hB3: lut_inv_sqrt = 16'h6231;
        8'hB4: lut_inv_sqrt = 16'h6214;
        8'hB5: lut_inv_sqrt = 16'h61F8;
        8'hB6: lut_inv_sqrt = 16'h61DB;
        8'hB7: lut_inv_sqrt = 16'h61BE;
        8'hB8: lut_inv_sqrt = 16'h61A2;
        8'hB9: lut_inv_sqrt = 16'h6186;
        8'hBA: lut_inv_sqrt = 16'h6169;
        8'hBB: lut_inv_sqrt = 16'h614D;
        8'hBC: lut_inv_sqrt = 16'h6131;
        8'hBD: lut_inv_sqrt = 16'h6115;
        8'hBE: lut_inv_sqrt = 16'h60F9;
        8'hBF: lut_inv_sqrt = 16'h60DD;
        8'hC0: lut_inv_sqrt = 16'h60C2;
        8'hC1: lut_inv_sqrt = 16'h60A6;
        8'hC2: lut_inv_sqrt = 16'h608B;
        8'hC3: lut_inv_sqrt = 16'h606F;
        8'hC4: lut_inv_sqrt = 16'h6054;
        8'hC5: lut_inv_sqrt = 16'h6039;
        8'hC6: lut_inv_sqrt = 16'h601E;
        8'hC7: lut_inv_sqrt = 16'h6003;
        8'hC8: lut_inv_sqrt = 16'h5FE8;
        8'hC9: lut_inv_sqrt = 16'h5FCD;
        8'hCA: lut_inv_sqrt = 16'h5FB2;
        8'hCB: lut_inv_sqrt = 16'h5F97;
        8'hCC: lut_inv_sqrt = 16'h5F7D;
        8'hCD: lut_inv_sqrt = 16'h5F62;
        8'hCE: lut_inv_sqrt = 16'h5F48;
        8'hCF: lut_inv_sqrt = 16'h5F2D;
        8'hD0: lut_inv_sqrt = 16'h5F13;
        8'hD1: lut_inv_sqrt = 16'h5EF9;
        8'hD2: lut_inv_sqrt = 16'h5EDF;
        8'hD3: lut_inv_sqrt = 16'h5EC5;
        8'hD4: lut_inv_sqrt = 16'h5EAB;
        8'hD5: lut_inv_sqrt = 16'h5E91;
        8'hD6: lut_inv_sqrt = 16'h5E77;
        8'hD7: lut_inv_sqrt = 16'h5E5D;
        8'hD8: lut_inv_sqrt = 16'h5E44;
        8'hD9: lut_inv_sqrt = 16'h5E2A;
        8'hDA: lut_inv_sqrt = 16'h5E11;
        8'hDB: lut_inv_sqrt = 16'h5DF7;
        8'hDC: lut_inv_sqrt = 16'h5DDE;
        8'hDD: lut_inv_sqrt = 16'h5DC5;
        8'hDE: lut_inv_sqrt = 16'h5DAC;
        8'hDF: lut_inv_sqrt = 16'h5D93;
        8'hE0: lut_inv_sqrt = 16'h5D7A;
        8'hE1: lut_inv_sqrt = 16'h5D61;
        8'hE2: lut_inv_sqrt = 16'h5D48;
        8'hE3: lut_inv_sqrt = 16'h5D2F;
        8'hE4: lut_inv_sqrt = 16'h5D17;
        8'hE5: lut_inv_sqrt = 16'h5CFE;
        8'hE6: lut_inv_sqrt = 16'h5CE6;
        8'hE7: lut_inv_sqrt = 16'h5CCD;
        8'hE8: lut_inv_sqrt = 16'h5CB5;
        8'hE9: lut_inv_sqrt = 16'h5C9D;
        8'hEA: lut_inv_sqrt = 16'h5C84;
        8'hEB: lut_inv_sqrt = 16'h5C6C;
        8'hEC: lut_inv_sqrt = 16'h5C54;
        8'hED: lut_inv_sqrt = 16'h5C3C;
        8'hEE: lut_inv_sqrt = 16'h5C24;
        8'hEF: lut_inv_sqrt = 16'h5C0C;
        8'hF0: lut_inv_sqrt = 16'h5BF5;
        8'hF1: lut_inv_sqrt = 16'h5BDD;
        8'hF2: lut_inv_sqrt = 16'h5BC5;
        8'hF3: lut_inv_sqrt = 16'h5BAE;
        8'hF4: lut_inv_sqrt = 16'h5B96;
        8'hF5: lut_inv_sqrt = 16'h5B7F;
        8'hF6: lut_inv_sqrt = 16'h5B68;
        8'hF7: lut_inv_sqrt = 16'h5B50;
        8'hF8: lut_inv_sqrt = 16'h5B39;
        8'hF9: lut_inv_sqrt = 16'h5B22;
        8'hFA: lut_inv_sqrt = 16'h5B0B;
        8'hFB: lut_inv_sqrt = 16'h5AF4;
        8'hFC: lut_inv_sqrt = 16'h5ADD;
        8'hFD: lut_inv_sqrt = 16'h5AC6;
        8'hFE: lut_inv_sqrt = 16'h5AAF;
        8'hFF: lut_inv_sqrt = 16'h5A99;
        default: lut_inv_sqrt = 16'h0000;
    endcase
endfunction
